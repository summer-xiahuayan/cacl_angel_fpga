`timescale 1ns/1ns
`include "cordic.v"
module cordic_angle_calc_tb ();

// ===================== �����ź� =====================
reg           clk;
reg           rst;
reg  signed [15:0] cx_in;
reg  signed [15:0] cy_in;

// ģ�����
wire signed [16:0] theta_1st_quad;  // ��һ���޽Ƕȣ����㣩
wire [1:0]         quadrant;        // ���ޱ��

// �ļ�����
integer cx_file, cy_file, out_file,true_angle_file;
integer read_cnt;
reg     file_end;

// ���Ƕȸ���
reg  signed [16:0] theta_1st_prev;
parameter EXT_NUM_ITERS = 19982;
real error [0:EXT_NUM_ITERS-1];
real error_sum=0.0;



// ===================== ʵ����ģ�� =====================
cordic_angle_calc u_angle_calc (
    .clk            (clk),
    .rst            (rst),
    .cx_in          (cx_in),
    .cy_in          (cy_in),
    .theta_1st_quad (theta_1st_quad),
    .quadrant       (quadrant)
);

// ===================== ʱ������ =====================
initial begin
    clk = 0;
    forever #5 clk = ~clk;  // 100MHz
end
real theta_1st_rad ;
real theta_1st_deg;
real true_angle;

        // �ڶ������������޼�����ʵ�Ƕȣ�������׶δ������򣡣�
real real_theta_rad;
real real_theta_deg;
// ===================== ���ģ���ӡ�����������ת��ʱ������ʵ�Ƕȣ� =====================
task print_result;
    input integer cnt;
    input signed [15:0] cx;
    input signed [15:0] cy;
    input [1:0] q;
    input signed [16:0] theta_1st;
    input real true_angle;
    real error_deg;
    begin
        // ��һ������һ���޽Ƕ�ת���㣨����ת����ʽ��
        theta_1st_rad = $itor(theta_1st) / 32768.0;
        theta_1st_deg = theta_1st_rad * 180.0 / 3.1415926535;

        // �ڶ������������޼�����ʵ�Ƕȣ�������׶δ������򣡣�      
        case (q)
            0: begin  // ��һ���ޣ�ֱ����
                real_theta_rad = theta_1st_rad;
                real_theta_deg = theta_1st_deg;
            end
            1: begin  // �ڶ����ޣ��� - ��һ���޽Ƕ�
                real_theta_rad = 3.1415926535/2 + theta_1st_rad;
                real_theta_deg = 180.0/2 + theta_1st_deg;
            end
            2: begin  // �������ޣ�-�� + ��һ���޽Ƕ�
                real_theta_rad = 3.1415926535 + theta_1st_rad;
                real_theta_deg = 180.0 + theta_1st_deg;
            end
            3: begin  // �������ޣ�-��һ���޽Ƕ�
                real_theta_rad = 3.1415926535*3/2+theta_1st_rad;
                real_theta_deg = 180.0*3/2+theta_1st_deg;
            end
        endcase
        error_deg= real_theta_deg-true_angle;
        // ��ӡ�����������ˣ�
        $display("���ݵ�%0d | cx=%0d, cy=%0d | ����%0d", cnt, cx, cy, q);
        $display("��һ���޽Ƕȣ�%f rad / %f ��", theta_1st_rad, theta_1st_deg);
        $display("FPGA����Ƕȣ�%f rad / %f ��", real_theta_rad, real_theta_deg);
        $display("MATLAB����Ƕȣ�%f ��", true_angle);
        $display("��%.6f ��\n", error_deg);
        error[cnt]=error_deg;
        error_sum=error_sum+error_deg;
        if (out_file != 0) begin
         $fwrite(out_file, "%f\n", real_theta_deg);
        end
        // д���ļ�����ѡ��
       // if (out_file != 0) begin
        //    $fwrite(out_file, "%d,%d,%d,%d,%f,%f\n", 
        //        cnt, cx, cy, q, real_theta_deg, true_angle);
       // end
    end
endtask

// ===================== ������ =====================
initial begin
    // ��ʼ��
    rst = 1;
    cx_in = 0;
    cy_in = 0;
    read_cnt = 0;
    file_end = 0;
    true_angle = 0;
    theta_1st_prev = 0;
    #20 rst = 0;

    // ���ļ�
    true_angle_file=$fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/angle_deg_360.txt", "r");
    cx_file  = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/cx_int16.txt", "r");
    cy_file  = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/cy_int16.txt", "r");
    out_file = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/angle_result.txt", "w");
    if (cx_file==0 || cy_file==0||true_angle_file==0) begin $display("�ļ���ʧ�ܣ�"); $stop; end
   // if (out_file!=0) $fwrite(out_file, "���ݵ�,cx,cy,����,FPGA����Ƕ�(rad),MATLAB����Ƕ�(��)\n");

    // ���ж�ȡ+���Ƕȸ���
    while (!file_end) begin
        @(posedge clk);
        
        // ��ȡ����
        if (!$feof(cx_file) && !$feof(cy_file)) begin
            $fscanf(cx_file, "%d", cx_in);
            $fscanf(cy_file, "%d", cy_in);
            read_cnt = read_cnt + 1;
        end else begin
            file_end = 1;
        end

        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        $fscanf(true_angle_file, "%f", true_angle);
        print_result(read_cnt, cx_in, cy_in, quadrant, theta_1st_quad,true_angle);
   
    end

    // ����
    $display("������ɣ�������%0d�����ݵ�", read_cnt);
    $display("ƽ����%.6f",error_sum/EXT_NUM_ITERS);
    $fclose(cx_file); $fclose(cy_file); $fclose(out_file);
    #100 $stop;
end

endmodule
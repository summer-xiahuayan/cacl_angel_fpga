// -----------------------------------------------------------------------------
// kf_angel_app_tb.v
// �������˲�Ӧ��ģ�飨kf_angel_app����ר�ò���ģ��
// ���ܣ�
//  1. ���ز������ݣ�measurements.txt/truth.txt��
//  2. ����kf_angel_appģ�飬ģ����ʵ��������
//  3. ��֤�˲������������������
// -----------------------------------------------------------------------------
`timescale 1ns/1ps

module kf_angel_app_tb();

  // =========================================================================
  // �������ã���Ӧ��ģ�鱣��һ�£�
  // =========================================================================
  parameter W          = 24;
  parameter FRAC       = 14;
  parameter NR         = 32;
  parameter ADDRW      = 5;
  parameter ROM_FILE   = "D:/DLS/LIBEROPRO/acc_filter/stimulus/kf_2d.mem";
  parameter TEST_ITERS = 5000;  // ���Ե������������޸ģ�

  // =========================================================================
  // �����źŶ���
  // =========================================================================
  // ʱ��/��λ
  reg              clk;
  reg              rst_n;
  // ģ������
  reg  [W-1:0]     meas_in;      // ģ�����ֵ����
  // ģ�����
  wire [W-1:0]     kf_pos_out;   // �˲���λ��
  wire [W-1:0]     kf_vel_out;   // �˲����ٶ�
  wire             data_out_valid;// �����Ч��־

  // �ڲ����Ա���
  real ext_meas [0:TEST_ITERS-1];  // ���صĲ���ֵ��ʵ����
  real ext_truth [0:TEST_ITERS-1]; // ���ص���ʵֵ��ʵ����
  real asic_pos  [0:TEST_ITERS-1]; // ģ�����λ�ã�ʵ����
  real asic_vel  [0:TEST_ITERS-1]; // ģ������ٶȣ�ʵ����
  integer iter;
  integer fd;
  integer cycle_count;

  // =========================================================================
  // ʵ��������ģ�飨kf_angel_app��
  // =========================================================================
  kf_angel_app #(
    .W(W),
    .FRAC(FRAC),
    .NR(NR),
    .ADDRW(ADDRW),
    .ROM_FILE(ROM_FILE)
  ) u_kf_angel_app (
    .clk(clk),
    .rst_n(rst_n),
    .meas_in(meas_in),
    .kf_pos_out(kf_pos_out),
    .kf_vel_out(kf_vel_out),
    .data_out_valid(data_out_valid)
  );

  // =========================================================================
  // ʱ�����ɣ�100MHz������5ns��
  // =========================================================================
  initial begin
    clk = 1'b0;
    forever #5 clk = ~clk;
  end

  // =========================================================================
  // �̶���?ʵ��ת�����������Ĺ��ߣ�
  // =========================================================================
  function [W-1:0] real_to_sm;
    input real x;
    reg sign;
    integer mag_int;
    begin
      sign = (x < 0.0);
      mag_int = (sign ? -x : x) * (1 << FRAC);
      real_to_sm = {sign, mag_int[W-2:0]};
    end
  endfunction

  function real sm_to_real;
    input [W-1:0] sm;
    real val;
    begin
      val = $itor(sm[W-2:0]) / (1 << FRAC);
      sm_to_real = sm[W-1] ? -val : val;
    end
  endfunction

 
  // =========================================================================
  // ������1�����ز������ݣ�measurements.txt / truth.txt��
  // =========================================================================
  task load_test_data;
    integer fd_meas, fd_truth;
    integer scan_ret;
    begin
      // ���ز���ֵ
      fd_meas = $fopen("D:/DLS/LIBEROPRO/acc_filter/stimulus/measurements.txt", "r");
      if (fd_meas == 0) begin
        $display("ERROR: �޷��� measurements.txt��");
        $finish;
      end
      for (iter = 0; iter < TEST_ITERS; iter = iter + 1) begin
        scan_ret = $fscanf(fd_meas, "%f", ext_meas[iter]);
      end
      $fclose(fd_meas);

      // ������ʵֵ
      fd_truth = $fopen("D:/DLS/LIBEROPRO/acc_filter/stimulus/kf_expected.txt", "r");
      if (fd_truth == 0) begin
        $display("ERROR: �޷��� truth.txt��");
        $finish;
      end
      for (iter = 0; iter < TEST_ITERS; iter = iter + 1) begin
        scan_ret = $fscanf(fd_truth, "%f %f", ext_truth[iter],asic_vel[iter]);
      end
      $fclose(fd_truth);

      $display("�ɹ����� %0d ��������ݣ�", TEST_ITERS);
    end
  endtask

  // =========================================================================
  // ������2����ӡ���Խ�������ͳ�ƣ�
  // =========================================================================
  task print_test_result;
    real sum_raw_err, sum_kf_err;
    real raw_mse, kf_mse;
    begin
      sum_raw_err = 0.0;
      sum_kf_err  = 0.0;

      // ���������MSE��
      for (iter = 0; iter < TEST_ITERS; iter = iter + 1) begin
        sum_raw_err = sum_raw_err + (ext_meas[iter] - ext_truth[iter])**2;
        sum_kf_err  = sum_kf_err  + (asic_pos[iter] - ext_truth[iter])**2;
      end
      raw_mse = sum_raw_err / TEST_ITERS;
      kf_mse  = sum_kf_err  / TEST_ITERS;

      // ��ӡͳ�ƽ��
      $display("\n==================== ���Խ��ͳ�� ====================");
      $display("ԭʼ����ֵ MSE��%.6f", raw_mse);
      $display("�˲���λ�� MSE��%.6f", kf_mse);
      $display("���������ʣ�%.1f%%", (1.0 - kf_mse/raw_mse)*100.0);
      $display("���һ�ε��������");
      $display("  �˲�λ�ã�%.6f | ��ʵλ�ã�%.6f | ��%.6f",
               asic_pos[TEST_ITERS-1], ext_truth[TEST_ITERS-1],
               abs(asic_pos[TEST_ITERS-1]-ext_truth[TEST_ITERS-1]));
      $display("  �˲��ٶȣ�%.6f", asic_vel[TEST_ITERS-1]);
    end
  endtask

  // =========================================================================
  // ������3������������ļ������ڻ�ͼ������
  // =========================================================================
  task export_result_to_file;
    begin
      fd = $fopen("D:/DLS/LIBEROPRO/acc_filter/stimulus/kf_app_test_result.txt", "w");
      if (fd == 0) begin
        $display("WARNING: �޷��������Խ���ļ���");
      //  return;
      end

      // д���ͷ
      $fwrite(fd, "Iter, Measured, Truth, KF_Pos, KF_Vel, Pos_Err\n");
      // д�����е������
      for (iter = 0; iter < TEST_ITERS; iter = iter + 1) begin
        $fwrite(fd, "%d,%.6f,%.6f,%.6f,%.6f,%.6f\n",
                iter+1, ext_meas[iter], ext_truth[iter],
                asic_pos[iter], asic_vel[iter],
                abs(asic_pos[iter]-ext_truth[iter]));
      end
      $fclose(fd);

      $display("\n���Խ���ѵ�������kf_app_test_result.txt");
    end
  endtask

  // =========================================================================
  // ��������������ֵ����
  // =========================================================================
  function real abs;
    input real x;
    begin
      abs = (x < 0) ? -x : x;
    end
  endfunction
 // =========================================================================
  // ����������
  // =========================================================================
  initial begin
    // --------------------------
    // 1. ��ʼ��
    // --------------------------
    $display("================================================================");
    $display("��ʼ���� kf_angel_app ģ�� - ����������%0d", TEST_ITERS);
    $display("================================================================");

    // ��λ�źų�ʼ��
    rst_n    = 1'b0;
    meas_in  = {W{1'b0}};
    cycle_count = 0;

    // ���ز������ݣ����ļ���ȡ��
    load_test_data();

    // --------------------------
    // 2. ��λ�ͷ�
    // --------------------------
    repeat(5) @(posedge clk);  // ��λ����5��ʱ��
    rst_n = 1'b1;
    $display("\n[�׶�1] ��λ�ͷţ�ģ������ʼ���׶�...");

    // --------------------------
    // 3. �ȴ�ģ���ʼ����ɣ�ǰ21��ʱ�ӣ�
    // --------------------------
    meas_in = real_to_sm(ext_meas[0]);
    repeat(21) @(posedge clk);
    $display("[�׶�2] ģ���ʼ����ɣ���ʼ�����������...");

    // --------------------------
    // 4. ѭ���������ֵ���ɼ����
    // --------------------------
    $display("\nIter |  �������ֵ  |  PYTHONֵ  |  �˲�λ��  |  λ�����  |  �˲��ٶ�");
    $display("-----|--------------|----------|------------|------------|----------");

    for (iter = 0; iter < TEST_ITERS; iter = iter + 1) begin
      // ���뵱ǰ����ֵ
      meas_in = real_to_sm(ext_meas[iter+1]);
      
      // �ȴ������Ч�����300��ʱ�ӳ�ʱ������
      cycle_count = 0;
      begin : wait_valid
        forever begin
          @(posedge clk);
          cycle_count = cycle_count + 1;
          
          // �����Ч���ɼ�����
          if (data_out_valid) begin
            asic_pos[iter] = sm_to_real(kf_pos_out);
            asic_vel[iter] = sm_to_real(kf_vel_out);
            
            // ��ӡ�ؼ����������ǰ10/��10/ÿ50�Σ�
            if (iter < 10 || iter >= TEST_ITERS-10 || (iter % 50 == 49)) begin
              $display("%4d |  %9.4f  | %8.4f |  %8.4f |  %8.6f | %8.4f",
                       iter+1, ext_meas[iter], ext_truth[iter],
                       asic_pos[iter], abs(asic_pos[iter]-ext_truth[iter]),
                       asic_vel[iter]);
            end
            disable wait_valid;
          end
          
          // ��ʱ����
          if (cycle_count > 300) begin
            $display("WARNING: ����%0d��ʱ��", iter);
            disable wait_valid;
          end
        end
      end
    end

    // --------------------------
    // 5. ���Խ��ͳ���뵼��
    // --------------------------
    print_test_result();
    export_result_to_file();

    // --------------------------
    // 6. ���Խ���
    // --------------------------
    $display("\n================================================================");
    $display("kf_angel_app ģ�������ɣ�");
    $display("================================================================");
    $finish;
  end

  // =========================================================================
  // ��ʱ���Ź�����ֹ��ѭ����
  // =========================================================================
  initial begin
    #(50_000_000);  // 50ms��ʱ
    $display("ERROR: ���Գ�ʱ��");
    $finish;
  end

endmodule
// -----------------------------------------------------------------------------
// pid_top_tb.v
// PID Controller ASIC Testbench (ƥ��ȫѭ��ָ���߼�)
// -----------------------------------------------------------------------------
`timescale 1ns/1ps

module pid_top_tb();

  // =========================================================================
  // Parameters (��ȫƥ�����PIDָ��ROM·��)
  // =========================================================================
  parameter ROM_FILE = "D:/DLS/LIBEROPRO/cacl_angel/stimulus/pid.mem";
  parameter EXT_NUM_ITERS = 19982;
  parameter W = 24;
  parameter FRAC = 14;
  parameter NR = 32;
  parameter ADDRW = 5;

  // =========================================================================
  // DUT Signals (����ԭ�ж���)
  // =========================================================================
  reg              clk;
  reg              rst_n;
  reg              START;
  reg  [W-1:0]     DATA_IN;
  reg  [ADDRW-1:0] DIR;
  reg              WRITE;
  wire             READY;
  wire [W-1:0]     DATA_OUT;
  reg              rom_we;
  reg  [7:0]       rom_waddr;
  reg  [15:0]      rom_wdata;
  reg  [7:0]       loop_addr;

  // Test data arrays (����PIDȫѭ���߼�)
  real ext_meas [0:EXT_NUM_ITERS-1];        // ����ֵ��ÿ��ѭ����ȡ��
  reg  [15:0]  ext_meas_int16 [0:EXT_NUM_ITERS-1]; // 16λ���Ͳ���ֵ
  real ext_setpoint [0:EXT_NUM_ITERS-1];    // ����ֵ��ÿ��ѭ����ȡ��
  // ASIC�������
  real asic_output [0:EXT_NUM_ITERS-1];     // PID���������(DB[8])
  reg  [23:0]  output_int16;
  reg  [15:0]  asic_output_int16 [0:EXT_NUM_ITERS-1];

  // PID���Ĳ�����ÿ��ѭ���������¼��ص�DB[0-2]��
  real Kp = 0.04;    // ����ϵ����1:1���ģ�
  real Ki = 0.01;   // ����ϵ��
  real Kd = 0;    // ΢��ϵ��

  // =========================================================================
  // DUT Instantiation (PIDģ��)
  // =========================================================================
`ifdef POST_SYN
  kf_top dut (
`else
  kf_top #(
    .W(W), .FRAC(FRAC), .NR(NR), .ADDRW(ADDRW), .ROM_FILE(ROM_FILE)
  ) dut (
`endif
    .clk(clk), .rst_n(rst_n), .START(START), .DATA_IN(DATA_IN),
    .DIR(DIR), .WRITE(WRITE), .READY(READY), .DATA_OUT(DATA_OUT),
    .rom_we(rom_we), .rom_waddr(rom_waddr), .rom_wdata(rom_wdata),
    .loop_addr(loop_addr)
  );

  // =========================================================================
  // Clock Generation (100 MHz)
  // =========================================================================
  initial clk = 0;
  always #5 clk = ~clk;

  // =========================================================================
  // Helper Functions (������ת��)
  // =========================================================================
  function [W-1:0] real_to_sm;
    input real x;
    reg sign;
    integer mag_int;
    begin
      sign = (x < 0.0);
      mag_int = (sign ? -x : x) * (1 << FRAC);
      real_to_sm = {sign, mag_int[W-2:0]};
    end
  endfunction

  function real sm_to_real;
    input [W-1:0] sm;
    real val;
    begin
      val = $itor(sm[W-2:0]) / (1 << FRAC);
      sm_to_real = sm[W-1] ? -val : val;
    end
  endfunction

  // =========================================================================
  // Extended PID Test - ��ȫƥ��ȫѭ��ָ���߼�
  // =========================================================================
  task test_ext_pid;
    integer iter, cycle_count, fd;
    integer scan_ret;
    real pid_output, error;
    real sum_err_sq, sum_output_sq;
    real y;
    begin
      // 3. ��ʼ��PID����������������ѭ���������ڼ��أ�
      loop_addr = 8'd2;  // LOOPָ������PC=0��ƥ�����ָ��PC=25: 0030��
      rst_n = 1;
      START = 1; @(posedge clk); START = 0; // ����ASIC

      // ��ʼ��ͳ�Ʊ���
      sum_err_sq = 0.0;
      sum_output_sq = 0.0;
      y = 0; // ��ʼ����ֵ���ɸ�����Ҫ������

      DATA_IN = real_to_sm(0.0);               @(posedge clk); // PC0: Load DB[0]=Kp
      DATA_IN = real_to_sm(0.0);               @(posedge clk); // PC1: Load DB[1]=Ki
      // 4. ���е�����ƥ��PIDȫѭ���߼���ÿ�ε���=1��PC0-25ѭ����
      for (iter = 0; iter < EXT_NUM_ITERS; iter = iter + 1) begin
        cycle_count = 0;
        // �����ڼ���PID������ƥ��ָ��PC0-4��Load�߼���
        DATA_IN = real_to_sm(Kp);               @(posedge clk); // PC0: Load DB[0]=Kp
        DATA_IN = real_to_sm(Ki);               @(posedge clk); // PC1: Load DB[1]=Ki
        DATA_IN = real_to_sm(Kd);               @(posedge clk); // PC2: Load DB[2]=Kd
        DATA_IN = real_to_sm(15.5);             @(posedge clk); // PC3: Load DB[3]=����ֵ
        DATA_IN = real_to_sm(y);                @(posedge clk); // PC4: Load DB[4]=����ֵ
        DATA_IN = 0; // ��������������

        // �ȴ�����PIDѭ����ɣ�PC����25: LOOPָ�
        begin : pid_loop_wait
          forever begin
            @(posedge clk);
            // ѭ��������־��PC=25�����LOOPָ��λ�ã�
            if (dut.Sequencer.pc == 8'd27) begin
              disable pid_loop_wait;
            end
            // ��ʱ����
            if (cycle_count > 300) begin 
              $display("WARNING: Timeout at iter %0d", iter);
              disable pid_loop_wait;
            end
          end
        end

        // ��ȡ����ѭ����PID�������ƥ������ڴ沼�֣�
        pid_output = sm_to_real(dut.Memory_Registers.Data_Bank_inst.mem[8]); // DB[8]=������
        y=4*pid_output+5;
        error      = sm_to_real(dut.Memory_Registers.Data_Bank_inst.mem[5]);  // DB[5]=��ǰ���
        output_int16 = dut.Memory_Registers.Data_Bank_inst.mem[8];
        

        // ��ӡ�ؼ��������
 
         $display("%4d | %8.2f ",iter + 1,pid_output);
      end

     
    end
  endtask

  // =========================================================================
  // Main Test (������)
  // =========================================================================
  initial begin
    $display("================================================================");
    $display("PID Controller ASIC Testbench (ƥ��ȫѭ��ָ���߼�)");
    $display("ָ��ѭ��: PC0(Load)��PC25(LOOP)��PC0 (����ѭ��)");
    $display("================================================================");

    // ��ʼ���ź�
    rst_n = 0; START = 0; DATA_IN = 0; DIR = 0; WRITE = 0;
    rom_we = 0; rom_waddr = 0; rom_wdata = 0; loop_addr = 0;

    // ��λ
    repeat(3) @(posedge clk);
    rst_n = 1;
    repeat(2) @(posedge clk);

    // ����PID��չ���ԣ�ƥ��ȫѭ���߼���
    test_ext_pid;

    $display("\n================================================================");
    $display("PID������� (ȫѭ���߼�ƥ��)");
    $display("================================================================\n");
    $finish;
  end

  // ��ʱ���Ź�
  initial begin
    #50000000;  // 50ms��ʱ����
    $display("ERROR: PID���Գ�ʱ!"); $finish;
  end

endmodule
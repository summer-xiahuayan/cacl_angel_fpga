`timescale 1ns/1ns
// ����ģ�飺cx/cy��һ�� + ȫ����ӳ�䵽��һ���� + ������ޱ��
module cordic_angle_calc (
    input           clk,            // ϵͳʱ��
    input           rst,            // ��λ������Ч��
    // ���룺16λ�з���cx/cyԭʼ����
    input  signed [15:0] cx_in,     // ��ӦMATLAB��cx_data
    input  signed [15:0] cy_in,     // ��ӦMATLAB��cy_data
    // �������һ���޽Ƕ� + ���ޱ��
    output signed [16:0] theta_1st_quad, // CORDIC����ĵ�һ���޽Ƕȣ�0~��/2��
    output reg [1:0]     quadrant        // ���ޱ�ţ�1=��һ��2=�ڶ���3=������4=���ģ�
);

// ===================== ��һ������������ =====================
// MATLAB��һ������
localparam signed [15:0] CX_DC        = 16'd17685;    // cxֱ������
localparam signed [15:0] CY_DC        = 16'd16800;    // cyֱ������
localparam signed [15:0] CX_NORM_COEFF= 16'd4990;     // cx��һ��ϵ��
localparam signed [15:0] CY_NORM_COEFF= 16'd5255;     // cy��һ��ϵ��
localparam DIV_SHIFT      = 10;                       // ��2^10 = ����10λ

// ===================== �ڶ�������һ�����㣨����ԭ���߼��� =====================
reg signed [15:0] cx_minus_dc;
reg signed [15:0] cy_minus_dc;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        cx_minus_dc <= 16'sd0;
        cy_minus_dc <= 16'sd0;
    end else begin
        cx_minus_dc <= cx_in - CX_DC;
        cy_minus_dc <= cy_in - CY_DC;
    end
end

reg signed [31:0] cx_mul_coeff;
reg signed [31:0] cy_mul_coeff;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        cx_mul_coeff <= 32'sd0;
        cy_mul_coeff <= 32'sd0;
    end else begin
        cx_mul_coeff <= cx_minus_dc * CX_NORM_COEFF;
        cy_mul_coeff <= cy_minus_dc * CY_NORM_COEFF;
    end
end

reg signed [16:0] cx_norm;
reg signed [16:0] cy_norm;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        cx_norm <= 17'sd0;
        cy_norm <= 17'sd0;
    end else begin
        cx_norm <= {cx_mul_coeff[31], cx_mul_coeff[25:10]} ;
        cy_norm <= {cy_mul_coeff[31], cy_mul_coeff[25:10]} ;
    end
end

// ===================== ����������ȷ�������ж� + ����ת��ӳ�䵽��һ���ޣ� =====================
reg [1:0] quadrant_comb;          // ����߼��ж�����
reg signed [16:0] cx_mapped;     // ӳ�䵽��һ���޵�cx
reg signed [16:0] cy_mapped;     // ӳ�䵽��һ���޵�cy

// ����߼��������ж� + ����ת�����ӳ٣�
always @(*) begin
    // Ĭ��ֵ�������ۺ���������
    quadrant_comb = 2'd1;
    cx_mapped = 17'sd0;
    cy_mapped = 17'sd0;

    // �ϸ����޹����ж� + ��׼����ת��ӳ�䵽��һ���ޣ�
    if (cx_norm >= 0 && cy_norm >= 0) begin
        // ��һ���ޣ�������ת��ֱ��ʹ��ԭ����
        quadrant_comb = 2'd0;
        cx_mapped = cx_norm;
        cy_mapped = cy_norm;
    end else if (cx_norm < 0 && cy_norm >= 0) begin
        // �ڶ����ޣ���ʱ��ת90�� �� (x,y) = (y, -x)
        quadrant_comb = 2'd1;
        cx_mapped = cy_norm;
        cy_mapped = -cx_norm;
    end else if (cx_norm < 0 && cy_norm < 0) begin
        // �������ޣ���ʱ��ת180�� �� (x,y) = (-x, -y)
        quadrant_comb = 2'd2;
        cx_mapped = -cx_norm;
        cy_mapped = -cy_norm;
    end else if (cx_norm >= 0 && cy_norm < 0) begin
        // �������ޣ���ʱ��ת270�� �� (x,y) = (-y, x)
        quadrant_comb = 2'd3;
        cx_mapped = -cy_norm;
        cy_mapped = cx_norm;
    end

    // ����0����ӳ���cx=0��ǿ����Ϊ1������CORDIC�����쳣��
    if (cx_mapped == 17'sd0) begin
        cx_mapped = 17'sd1;
    end
end

// ����ͬ��������߼�����Ĵ��������Ż�ʱ��
reg [1:0] quadrant_reg;
reg signed [16:0] cx_mapped_reg;
reg signed [16:0] cy_mapped_reg;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        quadrant <= 2'd0;
        cx_mapped_reg <= 17'sd0;
        cy_mapped_reg <= 17'sd0;
    end else begin
        quadrant <= quadrant_comb;
        cx_mapped_reg <= cx_mapped;
        cy_mapped_reg <= cy_mapped;
    end
end

// ===================== ���Ĳ���ʵ����CORDIC���������һ���޽Ƕȣ� =====================
cordic u_cordic (
    .clk      (clk),
    .rst      (rst),
    .x_i      (cx_mapped_reg),    // ӳ�䵽��һ���޵�cx
    .y_i      (cy_mapped_reg),    // ӳ�䵽��һ���޵�cy
    .theta_i  (17'sd0),           // VECTORģʽ�̶�Ϊ0
    .x_o      (),                 // ����
    .y_o      (),                 // ����
    .theta_o  (theta_1st_quad)    // �����һ���޽Ƕȣ�0~��/2��
);


endmodule
`timescale 1ns/1ns
module cordic_angle_calc_kf_tb ();

// ===================== �����ź� =====================
reg           clk;
reg           rst;
reg  signed [15:0] cx_in;
reg  signed [15:0] cy_in;

// ģ�����
wire signed [16:0] theta_1st_quad;  // ��һ���޽Ƕȣ����㣩
wire [1:0]         quadrant;        // ���ޱ��
wire               angle_valid;     // �����������Ч��־

// �ļ�����
integer cx_file, cy_file, out_file, true_angle_file;
integer read_cnt;
reg     file_end;

// ���ͳ��
parameter EXT_NUM_ITERS = 19982;
real error [0:EXT_NUM_ITERS-1];
real error_sum=0.0;

// ===================== ʵ����ģ�� =====================
cordic_angle_calc_kf u_angle_calc_kf (
    .clk            (clk),
    .rst            (rst),
    .cx_in          (cx_in),
    .cy_in          (cy_in),
    .theta_1st_quad (theta_1st_quad),
    .quadrant       (quadrant),
    .angle_valid    (angle_valid)
);

// ===================== ʱ������ =====================
initial begin
    clk = 0;
    forever #5 clk = ~clk;  // 100MHz������10ns��
end

// ===================== �Ƕ�ת�����ӡ���� =====================
real theta_1st_rad ;
real theta_1st_deg;
real true_angle;
real real_theta_rad;
real real_theta_deg;

// ��ӡ������񣨽�������Ч���ݣ�
task print_result;
    input integer cnt;
    input signed [15:0] cx;
    input signed [15:0] cy;
    input [1:0] q;
    input signed [16:0] theta_1st;
    input real true_angle;
    real error_deg;
    begin
        // ��һ���޽Ƕ�ת���㣨����ת����ʽ��
        theta_1st_rad = $itor(theta_1st) / 32768.0;
        theta_1st_deg = theta_1st_rad * 180.0 / 3.1415926535;

        // �������޼�����ʵ�Ƕ�
        case (q)
            0: begin  // ��һ���ޣ�ֱ����
                real_theta_rad = theta_1st_rad;
                real_theta_deg = theta_1st_deg;
            end
            1: begin  // �ڶ����ޣ���/2 + ��һ���޽Ƕ�
                real_theta_rad = 3.1415926535/2 + theta_1st_rad;
                real_theta_deg = 90.0 + theta_1st_deg;
            end
            2: begin  // �������ޣ��� + ��һ���޽Ƕ�
                real_theta_rad = 3.1415926535 + theta_1st_rad;
                real_theta_deg = 180.0 + theta_1st_deg;
            end
            3: begin  // �������ޣ�3��/2 + ��һ���޽Ƕ�
                real_theta_rad = 3.1415926535*3/2 + theta_1st_rad;
                real_theta_deg = 270.0 + theta_1st_deg;
            end
        endcase

        // ������
        error_deg = real_theta_deg - true_angle;
        error[cnt] = error_deg;
        error_sum = error_sum + error_deg;

        // ��ӡ���
        $display("=====================================");
        $display("���ݵ�%0d | �����Ч��YES", cnt);
        $display("cx=%0d, cy=%0d | ����%0d", cx, cy, q);
        $display("��һ���޽Ƕȣ�%f rad / %f ��", theta_1st_rad, theta_1st_deg);
        $display("FPGA(KF)����Ƕȣ�%f rad / %f ��", real_theta_rad, real_theta_deg);
        $display("MATLAB����Ƕȣ�%f ��", true_angle);
        $display("��%.6f ��", error_deg);
        $display("=====================================\n");

        // д���ļ�
        if (out_file != 0) begin
            $fwrite(out_file, "%d,%d,%d,%d,%f,%f\n", 
                cnt, cx, cy, q, real_theta_deg, true_angle);
        end
    end
endtask

// ===================== ���������̣����������������Чʱ�������룩 =====================
initial begin

    
    // ���ļ�
    true_angle_file = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/angle_filter_result.txt", "r");
    cx_file         = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/cx_int16.txt", "r");
    cy_file         = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/cy_int16.txt", "r");
    out_file        = $fopen("D:/DLS/LIBEROPRO/cacl_angel/stimulus/angle_result_kf.txt", "w");
    
    // �ļ��򿪼��
    if (cx_file==0 || cy_file==0 || true_angle_file==0) begin
        $display("�ļ���ʧ�ܣ�");
        $stop;
    end
    // д���ļ�ͷ
    if (out_file!=0) begin
        $fwrite(out_file, "���ݵ�,cx,cy,����,FPGA(KF)����Ƕ�(��),MATLAB����Ƕ�(��)\n");
    end

    // ��һ������ȡ��һ���ʼ����
    if (!$feof(cx_file) && !$feof(cy_file) && !$feof(true_angle_file)) begin
        $fscanf(cx_file, "%d", cx_in);
        $fscanf(cy_file, "%d", cy_in);
        $fscanf(true_angle_file, "%f", true_angle);
        read_cnt = read_cnt + 1;
    end else begin
        file_end = 1;
    end



    // ��ʼ��
    rst = 1;
  //  cx_in = 0;
   // cy_in = 0;
    read_cnt = 0;
    file_end = 0;
  //  true_angle = 0;
    repeat(5) @(posedge clk);  // ��λ����5��ʱ��
    rst = 0;
    // �����߼���ѭ���ȴ������Ч����Чʱ��ӡ+��������
    while (!file_end) begin
        // �ȴ�angle_valid��λ�������Ч��
      //  @(posedge clk iff angle_valid);
        @(posedge clk);
        if (angle_valid) begin
            
        // �����Чʱ����ӡ��ǰ���ݽ��
        print_result(read_cnt, cx_in, cy_in, quadrant, theta_1st_quad, true_angle);

        // �����Чʱ����ȡ��һ���������ݣ��������룩
        if (!$feof(cx_file) && !$feof(cy_file) && !$feof(true_angle_file)) begin
            $fscanf(cx_file, "%d", cx_in);
            $fscanf(cy_file, "%d", cy_in);
            $fscanf(true_angle_file, "%f", true_angle);
            read_cnt = read_cnt + 1;
        end else begin
            file_end = 1;  // �����ݿɶ�������ѭ��
        end
            
        end

    end

    // ���Խ�������
    $display("=====================================");
    $display("KF�汾������ɣ�������%0d����Ч���ݵ�", read_cnt-1);  // ��1����Ϊ���һ�ζ�ȡδ��ӡ
    $display("ƽ����%.6f ��", error_sum/(read_cnt-1));
    $display("=====================================");
    
    // �ر��ļ�
    $fclose(cx_file);
    $fclose(cy_file);
    $fclose(true_angle_file);
    $fclose(out_file);
    
    #100 $stop;
end

endmodule
// -----------------------------------------------------------------------------
// kf_angel_app.v
// �����������˲�Ӧ��ģ�飨����test_ext_kf�����߼���װ��
// ���ܣ�2D�������˲����̻���ʼ��ϵ���������Ⱪ¶ʱ��/��λ/����/����˿�
// ���룺ʱ�ӡ���λ������ֵ��24λ�̶��㣩
// ������˲���λ��/�ٶȣ�24λ�̶��㣩�������Ч��־
// -----------------------------------------------------------------------------
`timescale 1ns/1ps

module kf_angel_app
#(
  // �̶����������ԭ����ģ��һ�£�
  parameter W = 24,
  parameter FRAC = 14,
  parameter NR = 32,
  parameter ADDRW = 5,
  // ROM�ļ�·��������ʵ��·���޸ģ�
  parameter ROM_FILE = "D:/DLS/LIBEROPRO/acc_filter/stimulus/kf_2d.mem"
)
(
  input              clk,          // 100MHzʱ��
  input              rst_n,        // ����Ч��λ
  input  [W-1:0]     meas_in,      // �������ֵ��24λ�̶��㣬Q(23,14)��
  output reg [W-1:0] kf_pos_out,   // �˲���λ�������ͬ��ʽ��
  output reg [W-1:0] kf_vel_out,   // �˲����ٶ������ͬ��ʽ��
  output reg         data_out_valid// �����Ч��־���ߵ�ƽ��ʾ���ݿ��ã�
);

  // =========================================================================
  // �ڲ��źţ��Խ�ԭDUT�ӿڣ�
  // =========================================================================
  reg              START;
  reg  [W-1:0]     DATA_IN;
  reg  [ADDRW-1:0] DIR;
  reg              WRITE;
  wire             READY;
  wire [W-1:0]     DATA_OUT;
  wire             data_out_valid_dut; // DUT�����Ч
  reg  [7:0]       loop_addr;
  reg              rom_we;
  reg  [7:0]       rom_waddr;
  reg  [15:0]      rom_wdata;

  // ״̬���ƼĴ�������ʼ��/���У�
  reg [7:0]        init_cont;      // ��ʼ����������0~20��
  reg [15:0]       data_cont;      // �������������
  reg              init_done;      // ��ʼ����ɱ�־

  // =========================================================================
  // DUTʵ������ԭ�������˲�����ģ�飩
  // =========================================================================
  kf_angel_top #(
    .W(W), .FRAC(FRAC), .NR(NR), .ADDRW(ADDRW), .ROM_FILE(ROM_FILE)
  ) dut (
    .clk(clk), .rst_n(rst_n), .START(START), .DATA_IN(DATA_IN),
    .DIR(DIR), .WRITE(WRITE), .READY(READY), .DATA_OUT(DATA_OUT),
    .data_out_valid(data_out_valid_dut), .rom_we(rom_we), .rom_waddr(rom_waddr),
    .rom_wdata(rom_wdata), .loop_addr(loop_addr)
  );

  // =========================================================================
  // �̶���ת������������ԭ����ģ�飩
  // =========================================================================
  function [W-1:0] real_to_sm;
    input real x;
    reg sign;
    integer mag_int;
    begin
      sign = (x < 0.0);
      mag_int = (sign ? -x : x) * (1 << FRAC);
      real_to_sm = {sign, mag_int[W-2:0]};
    end
  endfunction

  // =========================================================================
  // ��ʼ���߼����̻�ϵ���������ⲿ���ã�
  // =========================================================================
  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      // ��λ��ʼ��
      START     <= 1'b0;
      DATA_IN   <= {W{1'b0}};
      loop_addr <= 8'd0;
      init_cont <= 8'd0;
      init_done <= 1'b0;
      rom_we    <= 1'b0;
      rom_waddr <= 8'd0;
      rom_wdata <= 16'd0;
      DIR       <= {ADDRW{1'b0}};
      WRITE     <= 1'b0;
    end else if (!init_done) begin
      // �׶�1�������ź�
      if (init_cont == 8'd0) begin
        loop_addr <= 8'd20;       // �̶�loop_addr=20��ԭ����ֵ��
        DATA_IN   <= real_to_sm(0.0);
        START     <= 1'b1;        // ����START
        init_cont <= init_cont + 1'b1;
      end
      // �׶�2����ʱ�Ӽ��ع̻���KF��ʼ��ϵ������21��������
      else begin
        START <= 1'b0;
        case(init_cont)
          8'd1:  DATA_IN <= real_to_sm(0.0);    // x1 ��ʼλ��
          8'd2:  DATA_IN <= real_to_sm(0.03);   // x2 ��ʼ�ٶ�
          8'd3:  DATA_IN <= real_to_sm(1.0);    // p11
          8'd4:  DATA_IN <= real_to_sm(0.0);    // p12
          8'd5:  DATA_IN <= real_to_sm(0.0);    // p21
          8'd6:  DATA_IN <= real_to_sm(1.0);    // p22
          8'd7:  DATA_IN <= real_to_sm(1.0);    // phi11
          8'd8:  DATA_IN <= real_to_sm(0.1);    // phi12
          8'd9:  DATA_IN <= real_to_sm(0.0);    // phi21
          8'd10: DATA_IN <= real_to_sm(1.0);    // phi22
          8'd11: DATA_IN <= real_to_sm(0.01);   // q11
          8'd12: DATA_IN <= real_to_sm(0.0);    // q12
          8'd13: DATA_IN <= real_to_sm(0.0);    // q21
          8'd14: DATA_IN <= real_to_sm(0.01);   // q22
          8'd15: DATA_IN <= real_to_sm(1.0);    // h1
          8'd16: DATA_IN <= real_to_sm(0.0);    // h2
          8'd17: DATA_IN <= real_to_sm(0.1);    // R
          8'd18: DATA_IN <= real_to_sm(0.0);    // g1
          8'd19: DATA_IN <= real_to_sm(0.0);    // g2
          8'd20: DATA_IN <= real_to_sm(0.0);    // u
          8'd21: begin
            DATA_IN  <= meas_in;   // ��һ������ֵ���ⲿ���룩
            init_done <= 1'b1;     // ��ʼ����ɣ��������н׶�
          end
          default: DATA_IN <= {W{1'b0}};
        endcase
        if (init_cont <= 8'd20) begin
          init_cont <= init_cont + 1'b1;
        end
      end
    end
  end

  // =========================================================================
  // ���н׶Σ���������/����߼�������ָ����ʱ��
  // =========================================================================
  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      kf_pos_out    <= {W{1'b0}};
      kf_vel_out    <= {W{1'b0}};
      data_out_valid<= 1'b0;
      data_cont     <= 16'd0;
      DATA_IN       <= {W{1'b0}};
    end else if (init_done) begin
      // ��ʼ����ɺ󣬰�data_out_valid_dut�������ݸ���
      if (data_out_valid_dut) begin
        // ����˲�������
        kf_pos_out    <= DATA_OUT;
        kf_vel_out    <= 'd0;//dut.Memory_Registers.Data_Bank_inst.mem[1]; // �ٶȴ��ڲ��洢��ȡ
        data_out_valid<= 1'b1;
        // ������һ������ֵ
        DATA_IN       <= meas_in;
        data_cont     <= data_cont + 1'b1;
      end else begin
        data_out_valid<= 1'b0;
      end
    end
  end

endmodule